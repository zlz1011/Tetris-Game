module pressed(ps2_key_pressed,ps2_out,sel,x1,y1,x2,y2,x3,y3,x4,y4);

	input ps2_key_pressed;
	input [7:0] ps2_out;
	input [2:0] sel;
	inout [5:0] x1,y1,x2,y2,x3,y3,x4,y4;
	
	
endmodule 